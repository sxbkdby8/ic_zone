module sync_clk_switch(
    input clk
);
endmodule