// module feedback_cdc(
//     input clk_src,
//     input clk_dst, 
//     input rst_n_src,
//     input rst_n_dst,
//     input din,
//     output dout
// )

//     wire 
//     gnrl_dffr #(1) src_sync_dffr1(din, data_sync1, clk_src, rst_n_src);

// endmodule